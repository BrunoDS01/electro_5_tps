module decode_latch(
	input wire [31:0] pc,
	input wire branch_prediction,
	input wire [4:0]  rs1,
	input wire [4:0]  rs2,
	input wire [4:0]  rd,
	input wire [9:0]  funct,
	input wire [31:0] imm,
	input wire [6:0]  opcode,

	input wire [2:0] instr_type,
	input wire save_to_reg,
	input wire rs1_used,
	input wire rs2_used,
	input wire immediate_used,
	input wire is_branch,
	input wire rd_memory,
	input wire wr_memory,

	
	input wire stg_clk,
	input wire stg_ena,
	input wire stg_x,
	input wire reset,
	
	output reg [31:0] pc_out,
	output reg branch_prediction_out,
	output reg [4:0]  rs1_out,
	output reg [4:0]  rs2_out,
	output reg [4:0]  rd_out,
	output reg [9:0]  funct_out,
	output reg [31:0] imm_out,
	output reg [6:0]  opcode_out,

	output reg [2:0] instr_type_out,
	
	output reg save_to_reg_out,
	output reg rs1_used_out,
	output reg rs2_used_out,
	output reg immediate_used_out,
	output reg is_branch_out,
	output reg rd_memory_out,
	output reg wr_memory_out
);

always @(posedge stg_clk or posedge reset) begin
	if(reset) begin
		pc_out <= 0;
		branch_prediction_out <= 0;
		rs1_out <= 0;
		rs2_out <= 0;
		rd_out <= 0;
		funct_out <= 0;
		imm_out <= 0;
		opcode_out <= 0;
		
		instr_type_out <= 0;
		
		save_to_reg_out <= 0;
		rs1_used_out <= 0;
		rs2_used_out <= 0;
		immediate_used_out <= 0;
		is_branch_out <= 0;
		rd_memory_out <= 0;
		wr_memory_out <= 0;
	end
	else begin
		pc_out <= pc;
		branch_prediction_out <= branch_prediction;
        rs1_out <= rs1;
        rs2_out <= rs2;
        rd_out <= rd;
        funct_out <= funct;
        imm_out <= imm;
        opcode_out <= opcode;

		  instr_type_out <= instr_type;
			
			
        save_to_reg_out <= save_to_reg;
        rs1_used_out <= rs1_used;
        rs2_used_out <= rs2_used;
        immediate_used_out <= immediate_used;
        is_branch_out <= is_branch;
        rd_memory_out <= rd_memory;
        wr_memory_out <= wr_memory;
	end
end

endmodule